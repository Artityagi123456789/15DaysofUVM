parameter WIDTH =16;
parameter DEPTH = 64;
parameter ADDR_WIDTH=$clog2(DEPTH);

class mem_common;
endclass
